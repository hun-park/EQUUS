module LUT (
    input   wire [19:00]    addr,
    output  reg  [39:00]    dout,
    output                  vital
);


always @(*) begin
    dout <= 40'd0;
    case(addr)
        20'd1 : dout <= {24'd102, 4'b0110, 4'b0000, 8'b00000000} ;
        20'd2 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd3 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd4 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd5 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd6 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd7 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd8 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd9 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd10 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd11 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd12 : dout <= {24'd63, 4'b0110, 4'b0000, 8'b00000000} ;
        20'd13 : dout <= {24'd95, 4'b0100, 4'b0000, 8'b00000000} ;
        20'd14 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd15 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd16 : dout <= {24'd63, 4'b0110, 4'b0000, 8'b00000000} ;
        20'd17 : dout <= {24'd95, 4'b0100, 4'b0000, 8'b00000000} ;
        20'd18 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd19 : dout <= {24'd47, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd20 : dout <= {24'd47, 4'b0000, 4'b0100, 8'b00010000} ;
        20'd21 : dout <= {24'd0, 4'b0010, 4'b0100, 8'b00100000} ;
        20'd22 : dout <= {24'd62, 4'b0010, 4'b0100, 8'b00010000} ;
        20'd23 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd24 : dout <= {24'd63, 4'b0110, 4'b0000, 8'b00000000} ;
        20'd25 : dout <= {24'd95, 4'b0100, 4'b0000, 8'b00000000} ;
        20'd26 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd27 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd28 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd29 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd30 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd31 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd32 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd33 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd34 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd35 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd36 : dout <= {24'd63, 4'b0110, 4'b0000, 8'b00000000} ;
        20'd37 : dout <= {24'd95, 4'b0100, 4'b0000, 8'b00000000} ;
        20'd38 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd39 : dout <= {24'd47, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd40 : dout <= {24'd47, 4'b0000, 4'b0100, 8'b00010000} ;
        20'd41 : dout <= {24'd0, 4'b0010, 4'b0100, 8'b00100000} ;
        20'd42 : dout <= {24'd62, 4'b0010, 4'b0100, 8'b00010000} ;
        20'd43 : dout <= {24'd95, 4'b0000, 4'b0000, 8'b00000000} ;
        20'd44 : dout <= {24'd63, 4'b0010, 4'b0000, 8'b00000000} ;
        20'd45 : dout <= {24'd0, 4'b0110, 4'b0000, 8'b00000000} ;
        20'd46 : dout <= {24'd82, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd47 : dout <= {24'd49, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd48 : dout <= {24'd50, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd49 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd50 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd51 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd52 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd53 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd54 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd55 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd56 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd57 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd58 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd59 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd60 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd61 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd62 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd63 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd64 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd65 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd66 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd67 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd68 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd69 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd70 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd71 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd72 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd73 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd74 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd75 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd76 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd77 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd78 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd79 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd80 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd81 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd82 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd83 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd84 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd85 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd86 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd87 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd88 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd89 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd90 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd91 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd92 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd93 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd94 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd95 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd96 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd97 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd98 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd99 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd100 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd101 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd102 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd103 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd104 : dout <= {24'd2, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd105 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd106 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd107 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd108 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd109 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd110 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd111 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd112 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd113 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd114 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd115 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd116 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd117 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd118 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd119 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd120 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd121 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd122 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd123 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd124 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd125 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd126 : dout <= {24'd37, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd127 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd128 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd129 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd130 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd131 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd132 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd133 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd134 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd135 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd136 : dout <= {24'd11, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd137 : dout <= {24'd3, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd138 : dout <= {24'd853, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd139 : dout <= {24'd3, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd140 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd141 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd142 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd143 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd144 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd145 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd146 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd147 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd148 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd149 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd150 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd151 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd152 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd153 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd154 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd155 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd156 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd157 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd158 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd159 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd160 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd161 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd162 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd163 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd164 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd165 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd166 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd167 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd168 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd169 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd170 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd171 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd172 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd173 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd174 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd175 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd176 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd177 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd178 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd179 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd180 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd181 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd182 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd183 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd184 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd185 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd186 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd187 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd188 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd189 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd190 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd191 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd192 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd193 : dout <= {24'd31, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd194 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd195 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd196 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd197 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd198 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd199 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd200 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd201 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd202 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd203 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd204 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd205 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd206 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd207 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd208 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd209 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd210 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd211 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd212 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd213 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd214 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd215 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd216 : dout <= {24'd31, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd217 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd218 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd219 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd220 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd221 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd222 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd223 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd224 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd225 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd226 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd227 : dout <= {24'd37, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd228 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd229 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd230 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd231 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd232 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd233 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd234 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd235 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd236 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd237 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd238 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd239 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd240 : dout <= {24'd33, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd241 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd242 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd243 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd244 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd245 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd246 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd247 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd248 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd249 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd250 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd251 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd252 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd253 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd254 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd255 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd256 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd257 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd258 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd259 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd260 : dout <= {24'd68, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd261 : dout <= {24'd2, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd262 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd263 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd264 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd265 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd266 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd267 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd268 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd269 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd270 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd271 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd272 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd273 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd274 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd275 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd276 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd277 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd278 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd279 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd280 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd281 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd282 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd283 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd284 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd285 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd286 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd287 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd288 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd289 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd290 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd291 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd292 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd293 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd294 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd295 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd296 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd297 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd298 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd299 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd300 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd301 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd302 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd303 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd304 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd305 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd306 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd307 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd308 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd309 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd310 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd311 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd312 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd313 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd314 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd315 : dout <= {24'd31, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd316 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd317 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd318 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd319 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd320 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd321 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd322 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd323 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd324 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd325 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd326 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd327 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd328 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd329 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd330 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd331 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd332 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd333 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd334 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd335 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd336 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd337 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd338 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd339 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd340 : dout <= {24'd33, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd341 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd342 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd343 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd344 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd345 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd346 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd347 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd348 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd349 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd350 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd351 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd352 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd353 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd354 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd355 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd356 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd357 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd358 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd359 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd360 : dout <= {24'd68, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd361 : dout <= {24'd2, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd362 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd363 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd364 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd365 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd366 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd367 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd368 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd369 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd370 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd371 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd372 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd373 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd374 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd375 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd376 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd377 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd378 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd379 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd380 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd381 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd382 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd383 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd384 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd385 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd386 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd387 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd388 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd389 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd390 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd391 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd392 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd393 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd394 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd395 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd396 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd397 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd398 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd399 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd400 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd401 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd402 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd403 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd404 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd405 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd406 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd407 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd408 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd409 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd410 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd411 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd412 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd413 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd414 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd415 : dout <= {24'd31, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd416 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd417 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd418 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd419 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd420 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd421 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd422 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd423 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd424 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd425 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd426 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd427 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd428 : dout <= {24'd35, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd429 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd430 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd431 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd432 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd433 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd434 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd435 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd436 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd437 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd438 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd439 : dout <= {24'd2, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd440 : dout <= {24'd34, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd441 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd442 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd443 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd444 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd445 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd446 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd447 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd448 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd449 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd450 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd451 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd452 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd453 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd454 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd455 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd456 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd457 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd458 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd459 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd460 : dout <= {24'd68, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd461 : dout <= {24'd2, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd462 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd463 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd464 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd465 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd466 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd467 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd468 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd469 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd470 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd471 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd472 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd473 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd474 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd475 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd476 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd477 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd478 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd479 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd480 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd481 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd482 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd483 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd484 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd485 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd486 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd487 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd488 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd489 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd490 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd491 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd492 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd493 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd494 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd495 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd496 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd497 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd498 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd499 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd500 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd501 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd502 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd503 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd504 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd505 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd506 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd507 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd508 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd509 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd510 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd511 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd512 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd513 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd514 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd515 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd516 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd517 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd518 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd519 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd520 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd521 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd522 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd523 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd524 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd525 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd526 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd527 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd528 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd529 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd530 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd531 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd532 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd533 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd534 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd535 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd536 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd537 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd538 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd539 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd540 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd541 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd542 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd543 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd544 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd545 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd546 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd547 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd548 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd549 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd550 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd551 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd552 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd553 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd554 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd555 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd556 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd557 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd558 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd559 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd560 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd561 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd562 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd563 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd564 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd565 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd566 : dout <= {24'd65535, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd567 : dout <= {24'd63892, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd568 : dout <= {24'd2, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd569 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd570 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd571 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd572 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd573 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd574 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd575 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd576 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd577 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd578 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd579 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd580 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd581 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd582 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd583 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd584 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd585 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd586 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd587 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd588 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd589 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd590 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd591 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd592 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd593 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd594 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd595 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd596 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd597 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd598 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd599 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd600 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd601 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd602 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd603 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd604 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd605 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd606 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd607 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd608 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd609 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd610 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd611 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd612 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd613 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd614 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd615 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd616 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd617 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd618 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd619 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd620 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd621 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd622 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd623 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd624 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd625 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd626 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd627 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd628 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd629 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd630 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd631 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd632 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd633 : dout <= {24'd2, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd634 : dout <= {24'd34, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd635 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd636 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd637 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd638 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd639 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd640 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd641 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd642 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd643 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd644 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd645 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd646 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd647 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd648 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd649 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd650 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd651 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd652 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd653 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd654 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd655 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd656 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd657 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd658 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd659 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd660 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd661 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd662 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd663 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd664 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd665 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd666 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd667 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd668 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd669 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd670 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd671 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd672 : dout <= {24'd33, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd673 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd674 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd675 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd676 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd677 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd678 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd679 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd680 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd681 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd682 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd683 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd684 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd685 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd686 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd687 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd688 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd689 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd690 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd691 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd692 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd693 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd694 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd695 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd696 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd697 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd698 : dout <= {24'd27, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd699 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd700 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd701 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd702 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd703 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd704 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd705 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd706 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd707 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd708 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd709 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd710 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd711 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd712 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd713 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd714 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd715 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd716 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd717 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd718 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd719 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd720 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd721 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd722 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd723 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd724 : dout <= {24'd34, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd725 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd726 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd727 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd728 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd729 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd730 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd731 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd732 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd733 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd734 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd735 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd736 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd737 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd738 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd739 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd740 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd741 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd742 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd743 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd744 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd745 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd746 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd747 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd748 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd749 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd750 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd751 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd752 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd753 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd754 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd755 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd756 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd757 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd758 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd759 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd760 : dout <= {24'd14, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd761 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd762 : dout <= {24'd21, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd763 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd764 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd765 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd766 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd767 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd768 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd769 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd770 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd771 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd772 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd773 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd774 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd775 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd776 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd777 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd778 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd779 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd780 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd781 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd782 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd783 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd784 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd785 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd786 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd787 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd788 : dout <= {24'd3360, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd789 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd790 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd791 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd792 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd793 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd794 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd795 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd796 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd797 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd798 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd799 : dout <= {24'd37, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd800 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd801 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd802 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd803 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd804 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd805 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd806 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd807 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd808 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd809 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd810 : dout <= {24'd19, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd811 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd812 : dout <= {24'd16, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd813 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd814 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd815 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd816 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd817 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd818 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd819 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd820 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd821 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd822 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd823 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd824 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd825 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd826 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd827 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd828 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd829 : dout <= {24'd10, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd830 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd831 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd832 : dout <= {24'd33345, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd833 : dout <= {24'd33345, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd834 : dout <= {24'd33345, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd835 : dout <= {24'd33345, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd836 : dout <= {24'd33345, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd837 : dout <= {24'd33345, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd838 : dout <= {24'd33345, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd839 : dout <= {24'd33345, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd840 : dout <= {24'd3, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd841 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd842 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd843 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd844 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd845 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd846 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd847 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd848 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd849 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd850 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd851 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd852 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd853 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd854 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd855 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd856 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd857 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd858 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd859 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd860 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd861 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd862 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd863 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd864 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd865 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd866 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd867 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd868 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd869 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd870 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd871 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd872 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd873 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd874 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd875 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd876 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd877 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd878 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd879 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd880 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd881 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd882 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd883 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd884 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd885 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd886 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd887 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd888 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd889 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd890 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd891 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd892 : dout <= {24'd37, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd893 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd894 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd895 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd896 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd897 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd898 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd899 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd900 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd901 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd902 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd903 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd904 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd905 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd906 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd907 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd908 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd909 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd910 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd911 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd912 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd913 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd914 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd915 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd916 : dout <= {24'd2, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd917 : dout <= {24'd34, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd918 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd919 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd920 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd921 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd922 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd923 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd924 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd925 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd926 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd927 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd928 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd929 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd930 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd931 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd932 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd933 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd934 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd935 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd936 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd937 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd938 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd939 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd940 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd941 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd942 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd943 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd944 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd945 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd946 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd947 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd948 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd949 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd950 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd951 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd952 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd953 : dout <= {24'd37, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd954 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd955 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd956 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd957 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd958 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd959 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd960 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd961 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd962 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd963 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd964 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd965 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd966 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd967 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd968 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd969 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd970 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd971 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd972 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd973 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd974 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd975 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd976 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd977 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd978 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd979 : dout <= {24'd27, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd980 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd981 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd982 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd983 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd984 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd985 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd986 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd987 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd988 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd989 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd990 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd991 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd992 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd993 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd994 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd995 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd996 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd997 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd998 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd999 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1000 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd1001 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1002 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1003 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1004 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1005 : dout <= {24'd34, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1006 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1007 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1008 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1009 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1010 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1011 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1012 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1013 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd1014 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1015 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1016 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1017 : dout <= {24'd36, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1018 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1019 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1020 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1021 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1022 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1023 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1024 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1025 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd1026 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1027 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1028 : dout <= {24'd3, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1029 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1030 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1031 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1032 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1033 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1034 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1035 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1036 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1037 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1038 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd1039 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1040 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1041 : dout <= {24'd37, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1042 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1043 : dout <= {24'd2, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1044 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1045 : dout <= {24'd1, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1046 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1047 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1048 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1049 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd1050 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1051 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1052 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1053 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1054 : dout <= {24'd30, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1055 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1056 : dout <= {24'd4, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1057 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1058 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1059 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b01000000} ;
        20'd1060 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b11000000} ;
        20'd1061 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1062 : dout <= {24'd0, 4'b0111, 4'b1000, 8'b10000000} ;
        20'd1063 : dout <= {24'd0, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1064 : dout <= {24'd0, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1065 : dout <= {24'd5, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1066 : dout <= {24'd1, 4'b1111, 4'b0000, 8'b00000000} ;
        20'd1067 : dout <= {24'd3360, 4'b0111, 4'b0000, 8'b00000000} ;
        20'd1068 : dout <= {24'hffffff, 4'b0000, 4'b0000, 8'b01010101};
        default : dout <= {24'h0, 4'b0000, 4'b0000, 8'b01010101};
    endcase
end
assign vital = 1'b1;
endmodule
